
--------***ROM 16x16x8(Q no:53)***--------
-------coded by Jenson and Salahudheen----

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.std_logic_arith.all;
--------------------------------------
entity ROM16x16x8 is
  port(
    clk,read,cs:in std_logic;
    add:in std_logic_vector(15 downto 0);
    data:out std_logic_vector(0 to 7));
end ROM16x16x8;
--------------------------------------
architecture Operation of ROM16x16x8 is
  
  type rom is array (0 to 15,0 to 15) of std_logic_vector(0 to 7);
  signal r:rom:=((("00111110"),("11111111"),("10101010"),("01010101"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("11111111"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("11111111"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("11111111"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")),
                (("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000"),
                ("00000000"),("00000000"),("00000000"),("00000000")));
  begin
    process(clk,read,cs,add)
      begin
        data<=r(conv_integer(add(15 downto 8)),conv_integer(add(7 downto 0)));
   end process; 
end Operation;