library ieee;
library Jenson_Salah;

use Jenson_Salah.Arrays.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
---------------------------------
entity KMap is
  port(
    noterms:in integer;
    
    
    
end KMap;
