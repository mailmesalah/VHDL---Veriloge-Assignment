library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
---------------------------------
entity ms is
  port(j,k,pr,clk,clr:in std_logic;
  q,qbar:inout std_logic);
end;
----------------------------------
architecture Op of ms is
signal ss,rm,ybar,q:std_logic:='1';
signal sm,rs,y,qbar:std_logic:='0';
begin
  
  
end;