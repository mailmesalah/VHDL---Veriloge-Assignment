library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
package Extras is
 
  --one dimentional integer array
  type integera is array(0 to 9) of integer range 0 to 100;
           
end Extras;  