
--------***RAM 16x16x8(Q no:53)***--------
-------coded by Jenson and Salahudheen----

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.std_logic_arith.all;
--------------------------------------
entity RAM16x16x8 is
  port(
    clk,read,cs,write:in std_logic;
    add:in std_logic_vector(15 downto 0);
    data:inout std_logic_vector(0 to 7));
end RAM16x16x8;
--------------------------------------
architecture Operation of RAM16x16x8 is
  
  type ram is array (0 to 15,0 to 15) of std_logic_vector(0 to 7);
  
  begin
    process(clk,read,cs,add,write)
      variable r:ram:=((("00111110"),("11111111"),("10101010"),("01010101"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("11111111"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("11111111"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("11111111"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")),
            (("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000"),
            ("00000000"),("00000000"),("00000000"),("00000000")));
      begin
        if (write='1' and clk='1' and cs='1') then
          r(conv_integer(add(15 downto 8)),conv_integer(add(7 downto 0))):=data;
        elsif (read='1' and cs='1' and clk='1') then
          data<=r(conv_integer(add(15 downto 8)),conv_integer(add(7 downto 0)));
        end if;
   end process; 
end Operation;